//-------------------------------------------------------------------------------------------------
// Lynx: Lynx 48K/96K/96Kscorpion implementation by Kyp
// https://github.com/Kyp069/lynx
//-------------------------------------------------------------------------------------------------
module audio
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      reset,
	input  wire      tape,
	input  wire[5:0] dac,
	output wire      q
);
//-------------------------------------------------------------------------------------------------

wire[9:0] mix = { 2'b00, {6{tape}} } + { 2'b00, dac };

dac #(.MSBI(9)) Dac
(
	.clock(clock  ),
	.reset(reset  ),
	.d    (mix    ),
	.q    (q      )
);

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
